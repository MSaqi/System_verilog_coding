module uart (
  /*------------------------------------------------------------------------------
  --  Comon signals CLK and rst_n
  ------------------------------------------------------------------------------*/
  input  logic        rst_n       ,
  input  logic        clk         ,
  /*------------------------------------------------------------------------------
  ------------------------------------------------------------------------------*/
  /*------------------------------------------------------------------------------
  --  UART TX Module Signals
  ------------------------------------------------------------------------------*/
  input  logic [31:0] data_in     ,
  input  logic        start       ,
  output reg          tx          ,
  output reg          tx_done     ,
  /*------------------------------------------------------------------------------
  ------------------------------------------------------------------------------*/
  /*------------------------------------------------------------------------------
  --  UART RX Module Signals
  ------------------------------------------------------------------------------*/
  input  logic        rx          ,
  output logic        rx_done     ,
  output reg   [31:0] dat_out     ,
  output reg   [ 3:0] parity_error
  /*------------------------------------------------------------------------------
  ------------------------------------------------------------------------------*/
);

  uart_tx tx_i (
    .clk    (clk    ),
    .rst_n  (rst_n  ),
    .start  (start  ),
    .data_in(data_in),
    .tx     (tx     ),
    .tx_done(tx_done)
  );

  uart_rx rx_i (
    .clk         (clk         ),
    .rst_n       (rst_n       ),
    .rx_done     (rx_done     ),
    .data_out    (dat_out     ),
    .rx          (rx          ),
    .parity_error(parity_error)
  );

endmodule