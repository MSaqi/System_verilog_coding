package uart_pkg;
  /*------------------------------------------------------------------------------
  --  ENUM
  ------------------------------------------------------------------------------*/
  typedef enum reg [2:0]{
    IDLE   = 3'b000,
    START  = 3'b001,
    DATA   = 3'b010,
    PARITY = 3'b011,
    STOP   = 3'b100
  } e_fsm_state;

  `define HIGH 1
  `define LOW 0
  /*------------------------------------------------------------------------------
  ------------------------------------------------------------------------------*/
endpackage